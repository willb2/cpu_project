

module controls(opcode, regDst, regWrite, aluSrc, pcSrc, memRead, memWrite, memToReg, aluOp);
	input [4:0] opcode;
	output regDst, regWrite, aluSrc, pcSrc, memRead, memWrite, memToReg;
	output [3:0] aluOp;

	


	




endmodule