

module controls(aluOp, data1, data2, result, zero);
	input [3:0] aluOp
	input [31:0] data1, data2;
	output [31:0] result;
	output zero;

	


endmodule