

module program_counter(address1, address2, mux, addressOut);
	input mux;
	input [31:0] address1, address2;
	output [31:0] addressOut;

	


endmodule