

module data_memory(memRead, memWrite, address, dataIn, dataOut);
	input memRead, memWrite;
	input [31:0] address, dataIn;
	output [31:0] dataOut;

	


endmodule