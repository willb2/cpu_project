

module adder(data1, data2, result);
	input [31:0] data1, data2;
	output [31:0] result;


endmodule