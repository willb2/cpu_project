

module instr_memory(address, instruction);
	input [31:0] address;
	output [31:0] instruction;

	


endmodule