

module top();




endmodule