

module registers(readReg1, readReg2, writeReg, readData1, readData2, writeData);
	input [4:0] readReg1, readReg2, writeReg;
	input [31:0] writeData;
	output [31:0] readData1, readData2;

	


endmodule